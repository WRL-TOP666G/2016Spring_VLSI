* File: FA4.pex.netlist
* Created: Tue Jun  7 17:55:14 2016
* Program "Calibre xRC"
* Version "v2012.2_26.20"
* 
.include "FA4.pex.netlist.pex"
.subckt FA4  C0 S0 S1 A0 A1 VDD S2 S3 A2 A3 GND B0 B1 C4 B2 B3
* 
* B3	B3
* B2	B2
* C4	C4
* B1	B1
* B0	B0
* GND	GND
* A3	A3
* A2	A2
* S3	S3
* S2	S2
* VDD	VDD
* A1	A1
* A0	A0
* S1	S1
* S0	S0
* C0	C0
M0 N_noxref_12_M0_d N_4_M0_g N_GND_M0_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M1 N_noxref_13_M1_d N_5_M1_g N_GND_M1_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M2 N_71_M2_d N_18_M2_g N_GND_M2_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07 AD=7.5e-14
+ AS=2.45e-13 PD=3e-07 PS=1.48e-06
M3 N_72_M3_d N_19_M3_g N_GND_M3_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07 AD=7.5e-14
+ AS=2.45e-13 PD=3e-07 PS=1.48e-06
M4 N_S0_M4_d N_18_M4_g N_noxref_12_M4_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M5 N_S1_M5_d N_19_M5_g N_noxref_13_M5_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M6 N_42_M6_d N_C0_M6_g N_71_M6_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=7.5e-14 PD=1.48e-06 PS=3e-07
M7 N_43_M7_d N_2_M7_g N_72_M7_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=7.5e-14 PD=1.48e-06 PS=3e-07
M8 N_noxref_12_M8_d N_44_M8_g N_S0_M8_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M9 N_noxref_13_M9_d N_45_M9_g N_S1_M9_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M10 N_GND_M10_d N_C0_M10_g N_noxref_12_M10_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M11 N_GND_M11_d N_2_M11_g N_noxref_13_M11_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M12 N_GND_M12_d N_C0_M12_g N_44_M12_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M13 N_GND_M13_d N_2_M13_g N_45_M13_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M14 N_73_M14_d N_42_M14_g N_GND_M14_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06
M15 N_74_M15_d N_43_M15_g N_GND_M15_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06
M16 N_4_M16_d N_18_M16_g N_GND_M16_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M17 N_5_M17_d N_19_M17_g N_GND_M17_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M18 N_2_M18_d N_48_M18_g N_73_M18_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07
M19 N_3_M19_d N_49_M19_g N_74_M19_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07
M20 N_noxref_22_M20_d N_6_M20_g N_GND_M20_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M21 N_noxref_23_M21_d N_7_M21_g N_GND_M21_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M22 N_18_M22_d N_A0_M22_g N_noxref_22_M22_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M23 N_19_M23_d N_A1_M23_g N_noxref_23_M23_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M24 N_noxref_22_M24_d N_46_M24_g N_18_M24_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M25 N_noxref_23_M25_d N_47_M25_g N_19_M25_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M26 N_GND_M26_d N_B0_M26_g N_noxref_22_M26_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M27 N_GND_M27_d N_B1_M27_g N_noxref_23_M27_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M28 N_75_M28_d N_A0_M28_g N_GND_M28_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06
M29 N_76_M29_d N_A1_M29_g N_GND_M29_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06
M30 N_GND_M30_d N_B0_M30_g N_46_M30_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M31 N_GND_M31_d N_B1_M31_g N_47_M31_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M32 N_48_M32_d N_B0_M32_g N_75_M32_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07
M33 N_49_M33_d N_B1_M33_g N_76_M33_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07
M34 N_6_M34_d N_A0_M34_g N_GND_M34_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M35 N_7_M35_d N_A1_M35_g N_GND_M35_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M36 N_noxref_27_M36_d N_8_M36_g N_GND_M36_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M37 N_noxref_28_M37_d N_9_M37_g N_GND_M37_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M38 N_77_M38_d N_33_M38_g N_GND_M38_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06
M39 N_78_M39_d N_34_M39_g N_GND_M39_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06
M40 N_S2_M40_d N_33_M40_g N_noxref_27_M40_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M41 N_S3_M41_d N_34_M41_g N_noxref_28_M41_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M42 N_52_M42_d N_3_M42_g N_77_M42_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07
M43 N_53_M43_d N_3_M43_g N_78_M43_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07
M44 N_noxref_27_M44_d N_54_M44_g N_S2_M44_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M45 N_noxref_28_M45_d N_55_M45_g N_S3_M45_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M46 N_GND_M46_d N_3_M46_g N_noxref_27_M46_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M47 N_GND_M47_d N_3_M47_g N_noxref_28_M47_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M48 N_GND_M48_d N_3_M48_g N_54_M48_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M49 N_GND_M49_d N_3_M49_g N_55_M49_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M50 N_79_M50_d N_52_M50_g N_GND_M50_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06
M51 N_80_M51_d N_53_M51_g N_GND_M51_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06
M52 N_8_M52_d N_33_M52_g N_GND_M52_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M53 N_9_M53_d N_34_M53_g N_GND_M53_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M54 N_3_M54_d N_59_M54_g N_79_M54_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07
M55 N_C4_M55_d N_60_M55_g N_80_M55_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07
M56 N_noxref_37_M56_d N_10_M56_g N_GND_M56_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M57 N_noxref_38_M57_d N_11_M57_g N_GND_M57_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M58 N_33_M58_d N_A2_M58_g N_noxref_37_M58_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M59 N_34_M59_d N_A3_M59_g N_noxref_38_M59_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M60 N_noxref_37_M60_d N_57_M60_g N_33_M60_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M61 N_noxref_38_M61_d N_58_M61_g N_34_M61_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
M62 N_GND_M62_d N_B2_M62_g N_noxref_37_M62_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M63 N_GND_M63_d N_B3_M63_g N_noxref_38_M63_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M64 N_81_M64_d N_A2_M64_g N_GND_M64_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06
M65 N_82_M65_d N_A3_M65_g N_GND_M65_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06
M66 N_GND_M66_d N_B2_M66_g N_57_M66_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M67 N_GND_M67_d N_B3_M67_g N_58_M67_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
M68 N_59_M68_d N_B2_M68_g N_81_M68_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07
M69 N_60_M69_d N_B3_M69_g N_82_M69_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07
M70 N_10_M70_d N_A2_M70_g N_GND_M70_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M71 N_11_M71_d N_A3_M71_g N_GND_M71_s N_GND_M0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
M72 N_VDD_M72_d N_4_M72_g N_noxref_16_M72_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M73 N_VDD_M73_d N_5_M73_g N_noxref_17_M73_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M74 N_42_M74_d N_18_M74_g N_VDD_M74_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M75 N_43_M75_d N_19_M75_g N_VDD_M75_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M76 N_noxref_63_M76_d N_18_M76_g N_VDD_M76_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M77 N_noxref_64_M77_d N_19_M77_g N_VDD_M77_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M78 N_VDD_M78_d N_C0_M78_g N_42_M78_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M79 N_VDD_M79_d N_2_M79_g N_43_M79_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M80 N_S0_M80_d N_44_M80_g N_noxref_63_M80_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M81 N_S1_M81_d N_45_M81_g N_noxref_64_M81_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M82 N_noxref_16_M82_d N_C0_M82_g N_S0_M82_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M83 N_noxref_17_M83_d N_2_M83_g N_S1_M83_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M84 N_VDD_M84_d N_C0_M84_g N_44_M84_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M85 N_VDD_M85_d N_2_M85_g N_45_M85_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M86 N_2_M86_d N_42_M86_g N_VDD_M86_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M87 N_3_M87_d N_43_M87_g N_VDD_M87_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M88 N_4_M88_d N_18_M88_g N_VDD_M88_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M89 N_5_M89_d N_19_M89_g N_VDD_M89_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M90 N_VDD_M90_d N_48_M90_g N_2_M90_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M91 N_VDD_M91_d N_49_M91_g N_3_M91_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M92 N_VDD_M92_d N_6_M92_g N_noxref_24_M92_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M93 N_VDD_M93_d N_7_M93_g N_noxref_25_M93_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M94 N_noxref_65_M94_d N_A0_M94_g N_VDD_M94_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M95 N_noxref_66_M95_d N_A1_M95_g N_VDD_M95_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M96 N_18_M96_d N_46_M96_g N_noxref_65_M96_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M97 N_19_M97_d N_47_M97_g N_noxref_66_M97_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M98 N_noxref_24_M98_d N_B0_M98_g N_18_M98_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M99 N_noxref_25_M99_d N_B1_M99_g N_19_M99_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M100 N_48_M100_d N_A0_M100_g N_VDD_M100_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M101 N_49_M101_d N_A1_M101_g N_VDD_M101_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M102 N_VDD_M102_d N_B0_M102_g N_46_M102_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M103 N_VDD_M103_d N_B1_M103_g N_47_M103_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M104 N_VDD_M104_d N_B0_M104_g N_48_M104_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M105 N_VDD_M105_d N_B1_M105_g N_49_M105_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M106 N_6_M106_d N_A0_M106_g N_VDD_M106_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M107 N_7_M107_d N_A1_M107_g N_VDD_M107_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M108 N_VDD_M108_d N_8_M108_g N_noxref_31_M108_s N_VDD_M73_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M109 N_VDD_M109_d N_9_M109_g N_noxref_32_M109_s N_VDD_M72_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M110 N_52_M110_d N_33_M110_g N_VDD_M110_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M111 N_53_M111_d N_34_M111_g N_VDD_M111_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M112 N_noxref_67_M112_d N_33_M112_g N_VDD_M112_s N_VDD_M73_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M113 N_noxref_68_M113_d N_34_M113_g N_VDD_M113_s N_VDD_M72_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M114 N_VDD_M114_d N_3_M114_g N_52_M114_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M115 N_VDD_M115_d N_3_M115_g N_53_M115_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M116 N_S2_M116_d N_54_M116_g N_noxref_67_M116_s N_VDD_M73_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M117 N_S3_M117_d N_55_M117_g N_noxref_68_M117_s N_VDD_M72_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M118 N_noxref_31_M118_d N_3_M118_g N_S2_M118_s N_VDD_M73_b P_18 L=1.8e-07
+ W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M119 N_noxref_32_M119_d N_3_M119_g N_S3_M119_s N_VDD_M72_b P_18 L=1.8e-07
+ W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M120 N_VDD_M120_d N_3_M120_g N_54_M120_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M121 N_VDD_M121_d N_3_M121_g N_55_M121_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M122 N_3_M122_d N_52_M122_g N_VDD_M122_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M123 N_C4_M123_d N_53_M123_g N_VDD_M123_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M124 N_8_M124_d N_33_M124_g N_VDD_M124_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M125 N_9_M125_d N_34_M125_g N_VDD_M125_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M126 N_VDD_M126_d N_59_M126_g N_3_M126_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M127 N_VDD_M127_d N_60_M127_g N_C4_M127_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M128 N_VDD_M128_d N_10_M128_g N_noxref_39_M128_s N_VDD_M73_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M129 N_VDD_M129_d N_11_M129_g N_noxref_40_M129_s N_VDD_M72_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M130 N_noxref_69_M130_d N_A2_M130_g N_VDD_M130_s N_VDD_M73_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M131 N_noxref_70_M131_d N_A3_M131_g N_VDD_M131_s N_VDD_M72_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M132 N_33_M132_d N_57_M132_g N_noxref_69_M132_s N_VDD_M73_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M133 N_34_M133_d N_58_M133_g N_noxref_70_M133_s N_VDD_M72_b P_18 L=1.8e-07
+ W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
M134 N_noxref_39_M134_d N_B2_M134_g N_33_M134_s N_VDD_M73_b P_18 L=1.8e-07
+ W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M135 N_noxref_40_M135_d N_B3_M135_g N_34_M135_s N_VDD_M72_b P_18 L=1.8e-07
+ W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M136 N_59_M136_d N_A2_M136_g N_VDD_M136_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M137 N_60_M137_d N_A3_M137_g N_VDD_M137_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M138 N_VDD_M138_d N_B2_M138_g N_57_M138_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M139 N_VDD_M139_d N_B3_M139_g N_58_M139_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
M140 N_VDD_M140_d N_B2_M140_g N_59_M140_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M141 N_VDD_M141_d N_B3_M141_g N_60_M141_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M142 N_10_M142_d N_A2_M142_g N_VDD_M142_s N_VDD_M73_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
M143 N_11_M143_d N_A3_M143_g N_VDD_M143_s N_VDD_M72_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
*
.include "FA4.pex.netlist.FA4.pxi"
*
.ends
*
*




.GLOBAL GND VDD
VGND GND 0v DC 0v
VVDD VDD GND DC 1.8v
V1 A0 GND PULSE( 0V 1.8V 0u 0u 0u 1u 2u )
V2 B0 GND PULSE( 0V 1.8V 0u 0u 0u 2u 4u )
V3 A1 GND PULSE( 0V 1.8V 0u 0u 0u 4u 8u )
V4 B1 GND PULSE( 0V 1.8V 0u 0u 0u 8u 16u )
V5 A2 GND PULSE( 0V 1.8V 0u 0u 0u 16u 32u )
V6 B2 GND PULSE( 0V 1.8V 0u 0u 0u 32u 64u )
V7 A3 GND PULSE( 0V 1.8V 0u 0u 0u 64u 128u )
V8 B3 GND PULSE( 0V 1.8V 0u 0u 0u 128u 256u )
V9 C0 GND PULSE( 0V 1.8V 0u 0u 0u 0u 0u )

XFA4 C0 S0 S1 A0 A1 VDD S2 S3 A2 A3 GND B0 B1 C4 B2 B3FA4

.protect
.lib 'cic018.l' TT
.unprotect
.options post
.tran 0.01u 250u
.end
