* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT XOR Y A B GND VDD
** N=10 EP=5 IP=0 FDC=12
M0 2 1 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-12820 $Y=-2370 $D=0
M1 Y A 2 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-12130 $Y=-2370 $D=0
M2 2 6 Y GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-11440 $Y=-2370 $D=0
M3 GND B 2 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-10750 $Y=-2370 $D=0
M4 GND B 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-9290 $Y=-2370 $D=0
M5 1 A GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-8600 $Y=-2370 $D=0
M6 VDD 1 4 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-12820 $Y=755 $D=1
M7 7 A VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=-12130 $Y=755 $D=1
M8 Y 6 7 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=-11440 $Y=755 $D=1
M9 4 B Y VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-10750 $Y=755 $D=1
M10 VDD B 6 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-9290 $Y=755 $D=1
M11 1 A VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-8600 $Y=755 $D=1
.ENDS
***************************************
