* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT FA4 C0 S0 S1 A0 A1 VDD S2 S3 A2 A3 GND B0 B1 C4 B2 B3
** N=82 EP=16 IP=0 FDC=144
M0 12 4 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-7740 $Y=-2070 $D=0
M1 13 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-7730 $Y=7010 $D=0
M2 71 18 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=-7330 $Y=5440 $D=0
M3 72 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=-7320 $Y=14520 $D=0
M4 S0 18 12 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-7050 $Y=-2070 $D=0
M5 S1 19 13 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-7040 $Y=7010 $D=0
M6 42 C0 71 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=-6850 $Y=5440 $D=0
M7 43 2 72 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=-6840 $Y=14520 $D=0
M8 12 44 S0 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-6360 $Y=-2070 $D=0
M9 13 45 S1 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-6350 $Y=7010 $D=0
M10 GND C0 12 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-5670 $Y=-2070 $D=0
M11 GND 2 13 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-5660 $Y=7010 $D=0
M12 GND C0 44 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-4210 $Y=-2070 $D=0
M13 GND 2 45 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-4200 $Y=7010 $D=0
M14 73 42 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=-3895 $Y=5440 $D=0
M15 74 43 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=-3885 $Y=14520 $D=0
M16 4 18 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-3520 $Y=-2070 $D=0
M17 5 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-3510 $Y=7010 $D=0
M18 2 48 73 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=-3415 $Y=5440 $D=0
M19 3 49 74 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=-3405 $Y=14520 $D=0
M20 22 6 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-885 $Y=-2070 $D=0
M21 23 7 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-875 $Y=7010 $D=0
M22 18 A0 22 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-195 $Y=-2070 $D=0
M23 19 A1 23 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-185 $Y=7010 $D=0
M24 22 46 18 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=495 $Y=-2070 $D=0
M25 23 47 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=505 $Y=7010 $D=0
M26 GND B0 22 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=1185 $Y=-2070 $D=0
M27 GND B1 23 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=1195 $Y=7010 $D=0
M28 75 A0 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=2455 $Y=5440 $D=0
M29 76 A1 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=2465 $Y=14520 $D=0
M30 GND B0 46 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=2645 $Y=-2070 $D=0
M31 GND B1 47 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=2655 $Y=7010 $D=0
M32 48 B0 75 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=2935 $Y=5440 $D=0
M33 49 B1 76 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=2945 $Y=14520 $D=0
M34 6 A0 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=3335 $Y=-2070 $D=0
M35 7 A1 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=3345 $Y=7010 $D=0
M36 27 8 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=7535 $Y=7010 $D=0
M37 28 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=7565 $Y=-2070 $D=0
M38 77 33 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=7945 $Y=14520 $D=0
M39 78 34 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=7975 $Y=5440 $D=0
M40 S2 33 27 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=8225 $Y=7010 $D=0
M41 S3 34 28 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=8255 $Y=-2070 $D=0
M42 52 3 77 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=8425 $Y=14520 $D=0
M43 53 3 78 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=8455 $Y=5440 $D=0
M44 27 54 S2 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=8915 $Y=7010 $D=0
M45 28 55 S3 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=8945 $Y=-2070 $D=0
M46 GND 3 27 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=9605 $Y=7010 $D=0
M47 GND 3 28 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=9635 $Y=-2070 $D=0
M48 GND 3 54 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=11065 $Y=7010 $D=0
M49 GND 3 55 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=11095 $Y=-2070 $D=0
M50 79 52 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=11380 $Y=14520 $D=0
M51 80 53 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=11410 $Y=5440 $D=0
M52 8 33 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=11755 $Y=7010 $D=0
M53 9 34 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=11785 $Y=-2070 $D=0
M54 3 59 79 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=11860 $Y=14520 $D=0
M55 C4 60 80 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=11890 $Y=5440 $D=0
M56 37 10 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=14390 $Y=7010 $D=0
M57 38 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=14420 $Y=-2070 $D=0
M58 33 A2 37 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=15080 $Y=7010 $D=0
M59 34 A3 38 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=15110 $Y=-2070 $D=0
M60 37 57 33 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=15770 $Y=7010 $D=0
M61 38 58 34 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=15800 $Y=-2070 $D=0
M62 GND B2 37 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=16460 $Y=7010 $D=0
M63 GND B3 38 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=16490 $Y=-2070 $D=0
M64 81 A2 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=17730 $Y=14520 $D=0
M65 82 A3 GND GND N_18 L=1.8e-07 W=5e-07 AD=7.5e-14 AS=2.45e-13 PD=3e-07 PS=1.48e-06 $X=17760 $Y=5440 $D=0
M66 GND B2 57 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=17920 $Y=7010 $D=0
M67 GND B3 58 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=17950 $Y=-2070 $D=0
M68 59 B2 81 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=18210 $Y=14520 $D=0
M69 60 B3 82 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=7.5e-14 PD=1.48e-06 PS=3e-07 $X=18240 $Y=5440 $D=0
M70 10 A2 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=18610 $Y=7010 $D=0
M71 11 A3 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=18640 $Y=-2070 $D=0
M72 VDD 4 16 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-7740 $Y=1425 $D=1
M73 VDD 5 17 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-7730 $Y=10505 $D=1
M74 42 18 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-7415 $Y=3510 $D=1
M75 43 19 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-7405 $Y=12590 $D=1
M76 63 18 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=-7050 $Y=1425 $D=1
M77 64 19 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=-7040 $Y=10505 $D=1
M78 VDD C0 42 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-6725 $Y=3510 $D=1
M79 VDD 2 43 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-6715 $Y=12590 $D=1
M80 S0 44 63 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=-6360 $Y=1425 $D=1
M81 S1 45 64 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=-6350 $Y=10505 $D=1
M82 16 C0 S0 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-5670 $Y=1425 $D=1
M83 17 2 S1 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-5660 $Y=10505 $D=1
M84 VDD C0 44 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-4210 $Y=1425 $D=1
M85 VDD 2 45 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-4200 $Y=10505 $D=1
M86 2 42 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-3980 $Y=3510 $D=1
M87 3 43 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-3970 $Y=12590 $D=1
M88 4 18 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-3520 $Y=1425 $D=1
M89 5 19 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-3510 $Y=10505 $D=1
M90 VDD 48 2 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-3290 $Y=3510 $D=1
M91 VDD 49 3 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-3280 $Y=12590 $D=1
M92 VDD 6 24 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-885 $Y=1425 $D=1
M93 VDD 7 25 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-875 $Y=10505 $D=1
M94 65 A0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=-195 $Y=1425 $D=1
M95 66 A1 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=-185 $Y=10505 $D=1
M96 18 46 65 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=495 $Y=1425 $D=1
M97 19 47 66 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=505 $Y=10505 $D=1
M98 24 B0 18 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=1185 $Y=1425 $D=1
M99 25 B1 19 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=1195 $Y=10505 $D=1
M100 48 A0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=2370 $Y=3510 $D=1
M101 49 A1 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=2380 $Y=12590 $D=1
M102 VDD B0 46 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=2645 $Y=1425 $D=1
M103 VDD B1 47 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=2655 $Y=10505 $D=1
M104 VDD B0 48 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=3060 $Y=3510 $D=1
M105 VDD B1 49 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=3070 $Y=12590 $D=1
M106 6 A0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=3335 $Y=1425 $D=1
M107 7 A1 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=3345 $Y=10505 $D=1
M108 VDD 8 31 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=7535 $Y=10505 $D=1
M109 VDD 9 32 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=7565 $Y=1425 $D=1
M110 52 33 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=7860 $Y=12590 $D=1
M111 53 34 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=7890 $Y=3510 $D=1
M112 67 33 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=8225 $Y=10505 $D=1
M113 68 34 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=8255 $Y=1425 $D=1
M114 VDD 3 52 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=8550 $Y=12590 $D=1
M115 VDD 3 53 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=8580 $Y=3510 $D=1
M116 S2 54 67 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=8915 $Y=10505 $D=1
M117 S3 55 68 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=8945 $Y=1425 $D=1
M118 31 3 S2 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=9605 $Y=10505 $D=1
M119 32 3 S3 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=9635 $Y=1425 $D=1
M120 VDD 3 54 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=11065 $Y=10505 $D=1
M121 VDD 3 55 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=11095 $Y=1425 $D=1
M122 3 52 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=11295 $Y=12590 $D=1
M123 C4 53 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=11325 $Y=3510 $D=1
M124 8 33 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=11755 $Y=10505 $D=1
M125 9 34 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=11785 $Y=1425 $D=1
M126 VDD 59 3 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=11985 $Y=12590 $D=1
M127 VDD 60 C4 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=12015 $Y=3510 $D=1
M128 VDD 10 39 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=14390 $Y=10505 $D=1
M129 VDD 11 40 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=14420 $Y=1425 $D=1
M130 69 A2 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=15080 $Y=10505 $D=1
M131 70 A3 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=15110 $Y=1425 $D=1
M132 33 57 69 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=15770 $Y=10505 $D=1
M133 34 58 70 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=15800 $Y=1425 $D=1
M134 39 B2 33 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=16460 $Y=10505 $D=1
M135 40 B3 34 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=16490 $Y=1425 $D=1
M136 59 A2 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=17645 $Y=12590 $D=1
M137 60 A3 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=17675 $Y=3510 $D=1
M138 VDD B2 57 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=17920 $Y=10505 $D=1
M139 VDD B3 58 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=17950 $Y=1425 $D=1
M140 VDD B2 59 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=18335 $Y=12590 $D=1
M141 VDD B3 60 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=18365 $Y=3510 $D=1
M142 10 A2 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=18610 $Y=10505 $D=1
M143 11 A3 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=18640 $Y=1425 $D=1
.ENDS
***************************************
